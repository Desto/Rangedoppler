-- RDA highest level architecture